*****Single NMOS Transistor (Id-Vd) ***

*** circuit description ***


m1 2 1 0 0 nmos1 L=1u W=10u

vgs 1 0 0 
vds 2 0 0 

.control
run
dc vds 0 5 0.05 vgs 0 5 0.5 
plot i(vds)
.endc


* Basic Level 1 default model for nchan
.MODEL nmos1 NMOS

* Basic Level 1 default model for pchan
.MODEL pmos1 PMOS

* Level 2 model nchan model for CN20
.MODEL CMOSN NMOS LEVEL=2 PHI=0.600000 TOX=4.3500E-08 XJ=0.200000U TPG=1
+ VTO=0.8756 DELTA=8.5650E+00 LD=2.3950E-07 KP=4.5494E-05 
+ UO=573.1 UEXP=1.5920E-01 UCRIT=5.9160E+04 RSH=1.0310E+01 
+ GAMMA=0.4179 NSUB=3.3160E+15 NFS=8.1800E+12 VMAX=6.0280E+04 
+ LAMBDA=2.9330E-02 CGDO=2.8518E-10 CGSO=2.8518E-10 
+ CGBO=4.0921E-10 CJ=1.0375E-04 MJ=0.6604 CJSW=2.1694E-10 
+ MJSW=0.178543 PB=0.800000
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is -4.0460E-07

* Level 2 model pchan model for CN20
.MODEL CMOSP PMOS LEVEL=2 PHI=0.600000 TOX=4.3500E-08 XJ=0.200000U TPG=-1
+ VTO=-0.8889 DELTA=4.8720E+00 LD=2.9230E-07 KP=1.5035E-05 
+ UO=189.4 UEXP=2.7910E-01 UCRIT=9.5670E+04 RSH=1.8180E+01 
+ GAMMA=0.7327 NSUB=1.0190E+16 NFS=6.1500E+12 VMAX=9.9990E+05 
+ LAMBDA=4.2290E-02 CGDO=3.4805E-10 CGSO=3.4805E-10 
+ CGBO=4.0305E-10 CJ=3.2456E-04 MJ=0.6044 CJSW=2.5430E-10 
+ MJSW=0.244194 PB=0.800000
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is -3.6560E-07

* BSIM model for n-channel CN20
.MODEL CMOSNB NMOS LEVEL=4 
+VFB=-9.73820E-01, LVFB=3.67458E-01,WVFB=-4.72340E-02
+phi=7.46556E-01,lphi=-1.92454E-24, wphi=8.06093E-24
+k1=1.49134E+00,lk1=-4.98139E-01, wk1=2.78225E-01
+k2=3.15199E-01,lk2=-6.95350E-02,wk2=-1.40057E-01
+eta=-1.19300E-02, leta=5.44713E-02,weta=-2.67784E-02
+muz=5.98328E+02,dl=6.38067E-001,dw=1.35520E-001
+u0=5.27788E-02, lu0=4.85686E-02,wu0=-8.55329E-02
+u1=1.09730E-01, lu1=7.28376E-01,wu1=-4.22283E-01
+x2mz=7.18857E+00,lx2mz=-2.47335E+00, wx2mz=7.12327E+01
+x2e=-3.00000E-03,lx2e=-7.20276E-03,wx2e=-5.57093E-03
+x3e=3.71969E-04,lx3e=-3.16123E-03,wx3e=-3.80806E-03
+x2u0=1.30153E-03, lx2u0=3.81838E-04, wx2u0=2.53131E-02
+x2u1=-2.04836E-02, lx2u1=3.48053E-02, wx2u1=4.44747E-02
+mus=7.79064E+02, lmus=3.62270E+02,wmus=-2.71207E+02
+x2ms=-2.65485E+00, lx2ms=3.68637E+01, wx2ms=1.12899E+02
+x3ms=1.18139E+01, lx3ms=7.24951E+01,wx3ms=-5.25361E+01
+x3u1=2.12924E-02, lx3u1=5.85329E-02,wx3u1=-5.29634E-02
+tox=4.35000E-002, temp=2.70000E+01, vdd=5.00000E+00  
+cgdo=3.79886E-010,cgso=3.79886E-010,cgbo=3.78415E-010
+xpart=1.00000E+000
+n0=1.00000E+000 ln0=0.00000E+000 wn0=0.00000E+000 
+nb=0.00000E+000 lnb=0.00000E+000 wnb=0.00000E+000 
+nd=0.00000E+000 lnd=0.00000E+000 wnd=0.00000E+000 
+rsh=27.9    cj=1.037500e-04    cjsw=2.169400e-10  js=1.000000e-08    pb=0.8    
+pbsw=0.8    mj=0.66036    mjsw=0.178543    wdf=0    dell=0

* BSIM model for p-channel CN20
.MODEL CMOSPB PMOS LEVEL=4
+ vfb=-2.65334E-01, lvfb=6.50066E-02, wvfb=1.48093E-01
+ phi=6.75823E-01,lphi=-1.61406E-24, wphi=8.03764E-24
+ k1=5.68962E-01, lk1=3.88845E-02,wk1=-5.33948E-02
+ k2=-5.52938E-02, lk2=1.17906E-01,wk2=-6.89149E-02
+ eta=-1.51784E-02, leta=5.87976E-02,weta=-7.51570E-04
+ muz=2.10669E+02,dl=8.44240E-001,dw=1.62551E-001
+ u0=1.04713E-01, lu0=5.50950E-02,wu0=-7.56659E-02
+ u1=1.46638E-02, lu1=2.13581E-01,wu1=-1.22509E-01
+ x2mz=8.76354E+00,lx2mz=-3.64793E+00, wx2mz=4.30934E+00
+ x2e=-2.13631E-03,lx2e=-2.94140E-03,wx2e=-2.48293E-03
+ x3e=2.78813E-04,lx3e=-1.60711E-03,wx3e=-4.57237E-03
+ x2u0=3.93706E-03,lx2u0=-5.66051E-04, wx2u0=5.69621E-04
+ x2u1=1.07707E-04, lx2u1=8.85125E-03, wx2u1=1.71537E-03
+ mus=2.06464E+02, lmus=1.39151E+02,wmus=-4.95671E+01
+ x2ms=5.86401E+00, lx2ms=6.98887E+00, wx2ms=5.55782E+00
+ x3ms=-2.03430E-01, lx3ms=1.16170E+01,wx3ms=-3.44342E+00
+ x3u1=-1.17893E-02, lx3u1=5.72098E-04, wx3u1=8.29791E-03
+ tox=4.35000E-002, temp=2.70000E+01, vdd=5.00000E+00   
+ cgdo=5.02635E-010,cgso=5.02635E-010,cgbo=3.85017E-010
+ xpart=1.00000E+000
+ n0=1.00000E+000,ln0=0.00000E+000,wn0=0.00000E+000
+ nb=0.00000E+000,lnb=0.00000E+000,wnb=0.00000E+000
+ nd=0.00000E+000,lnd=0.00000E+000,wnd=0.00000E+000
+ rsh=54.7,    cj=3.245600e-04,    cjsw=2.543000e-10,    js=1.000000e-08,    pb=0.8
+ pbsw=0.8,    mj=0.60438,    mjsw=0.244194,    wdf=0,    dell=0


* Lateral BJT model for CN20
.MODEL BN2X1 NPN
+ BF=82 IS=1.588E-16 NF=9.9563E-01 NE=1.3356 VAF=57.1
+ IKF=2.3067E-02 ISE=1.267E-16 RE=12.7 RC=420.00 RB=1.213E+03
+ RBM=7.53 ISC=3.363E-15 NC=1.0202
+ CJE=0.1952E-12 MJE=0.5050 VJE=0.85 CJC=0.18815E-12 MJC=0.4990 VJC=0.80
+ CJS=0.2326E-12 MJS=0.2033 VJS=0.70

* Level 3 SPICE model for CMOS14TB 0.5 um
.MODEL CMOSN5 NMOS LEVEL=3 PHI=0.700000 
+ TOX=9.6000E-09 XJ=0.200000U TPG=1
+ VTO=0.7118 DELTA=2.3060E-01 LD=2.9830E-08 KP=1.8201E-04 
+ UO=506.0 THETA=1.9090E-01 RSH=1.8940E+01 GAMMA=0.6051 
+ NSUB=1.4270E+17 NFS=7.1500E+11 VMAX=2.4960E+05 ETA=2.5510E-02 
+ KAPPA=1.8530E-01 CGDO=9.0000E-11 CGSO=9.0000E-11 
+ CGBO=3.7295E-10 CJ=6.02E-04 MJ=0.805 CJSW=2.0E-11 
+ MJSW=0.761 PB=0.99
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is 3.5700E-07

* Level 4 (BSIM) SPICE model for CMOS14TB 0.5 um
.MODEL CMOSNB5 NMOS LEVEL=4 
+ vfb=-9.65360E-01   	lvfb= 4.11254E-02   	wvfb=-1.21737E-01
+ phi= 9.02436E-01   	lphi= 0.00000E+00   	wphi= 0.00000E+00
+ k1=  9.33674E-01  	lk1= -8.15872E-02   	wk1=  2.03526E-01
+ k2=  7.39228E-02   	lk2=  1.48295E-02   	wk2=  5.89097E-02
+ eta=-2.77969E-03   	leta= 1.12296E-02   	weta= 1.25263E-03
+ muz= 4.71133E+02   	dl=   1.57937E-001  	dw=   4.09563E-001
+ u0=  1.98427E-01  	lu0=  1.54850E-01   	wu0= -1.05429E-01
+ u1=  3.39403E-02   	lu1=  3.59469E-02  	wu1= -5.00497E-03
+ x2mz=1.25728E+01 	lx2mz=-1.24115E+01  	wx2mz=1.77657E+01
+ x2e=-9.95217E-05   	lx2e=-5.16949E-03   	wx2e= 2.83253E-03
+ x3e=-4.27269E-04   	lx3e=-1.62632E-03   	wx3e=-1.60797E-03
+ x2u0=-9.02747E-04  	lx2u0=-1.66946E-02  	wx2u0=2.48458E-02
+ x2u1=-7.29822E-04  	lx2u1=2.38803E-03   	wx2u1=-9.76918E-04
+ mus=5.36631E+02    	lmus=2.18647E+01    	wmus=4.43373E+00
+ x2ms=5.97403E+00 	lx2ms=-7.67105E+00  	wx2ms=2.19614E+01
+ x3ms=7.60054E+00 	lx3ms=4.73779E+00   	wx3ms=2.59952E+00
+ x3u1=1.75532E-02   	lx3u1=-1.21628E-03  	wx3u1=-5.95548E-04
+ tox=9.60000E-003   	temp=2.70000E+01    	vdd=3.30000E+00
+ cgdo=4.26077E-010  	cgso=4.26077E-010   	cgbo=4.01709E-010
+ xpart=1.00000E+000
+ n0=1.00000E+000    	ln0=0.00000E+000    	wn0=0.00000E+000
+ nb=0.00000E+000    	lnb=0.00000E+000    	wnb=0.00000E+000
+ nd=0.00000E+000    	lnd=0.00000E+000    	wnd=0.00000E+000
+ rsh=2    cj=6.02e-04    cjsw=2.0e-11    js=1e-08  pb=0.99
+ pbsw=0.99    mj=0.805    mjsw=0.761    wdf=0    dell=0

* Level 3 SPICE model for CMOS14TB 0.5 um
.MODEL CMOSP5 PMOS LEVEL=3 PHI=0.700000 
+ TOX=9.6000E-09 XJ=0.200000U TPG=-1
+ VTO=-0.9016 DELTA=4.2020E-01 LD=4.3860E-08 KP=4.1582E-05 
+ UO=115.6 THETA=3.7990E-02 RSH=9.0910E-02 GAMMA=0.4496 
+ NSUB=7.8780E+16 NFS=6.4990E+11 VMAX=2.3130E+05 ETA=2.8580E-02 
+ KAPPA=9.9270E+00 CGDO=9.0000E-11 CGSO=9.0000E-11 
+ CGBO=3.6835E-10 CJ=9.34E-04 MJ=0.491 CJSW=2.41E-10 
+ MJSW=0.222 PB=0.90
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is 3.4860E-07

* Level 4 (BSIM) SPICE model for CMOS14TB 0.5 um
.MODEL CMOSPB5 PMOS LEVEL=4
+ vfb=-2.80568E-01   	lvfb=5.70163E-02    	wvfb=-6.17493E-02
+ phi=8.14689E-01    	lphi=0.00000E+00    	wphi=0.00000E+00
+ k1=4.52973E-01     	lk1=-9.19899E-02    	wk1=1.20834E-01
+ k2=-9.42157E-03    	lk2=-2.25562E-03    	wk2=3.13315E-02
+ eta=-7.03956E-03  	leta=1.92833E-02    	weta=5.45445E-05
+ muz=1.36047E+02    	dl=1.85988E-001     	dw=4.32366E-001
+ u0=1.93813E-01     	lu0=6.02231E-02     	wu0=-4.90734E-02
+ u1=8.52399E-03     	lu1=2.60545E-02     	wu1=-6.34371E-03
+ x2mz=7.96258E+00 	lx2mz=-2.15761E+00  	wx2mz=2.30663E+00
+ x2e=4.37912E-04    	lx2e=-1.60046E-03   	wx2e=-3.86750E-04
+ x3e=-3.52725E-04   	lx3e=-4.09096E-04   	wx3e=-2.53471E-03
+ x2u0=1.18873E-02   	lx2u0=-4.81760E-03  	wx2u0=8.80040E-03
+ x2u1=2.26591E-03   	lx2u1=7.96828E-04   	wx2u1=-4.70527E-04
+ mus=1.44421E+02    	lmus=1.63665E+01    	wmus=-7.31189E-01
+ x2ms=8.18970E+00 	lx2ms=-1.25158E+00  	wx2ms=3.62233E+00
+ x3ms=7.29640E-01  	lx3ms=1.15206E+00   	wx3ms=1.02833E+00
+ x3u1=-3.51521E-03  	lx3u1=-3.12374E-03  	wx3u1=3.48134E-03
+ tox=9.60000E-003   	temp=2.70000E+01    	vdd=3.30000E+00
+ cgdo=5.01753E-010  	cgso=5.01753E-010   	cgbo=4.14187E-010
+ xpart=1.00000E+000  
+ n0=1.00000E+000    	ln0=0.00000E+000    	wn0=0.00000E+000
+ nb=0.00000E+000    	lnb=0.00000E+000    	wnb=0.00000E+000
+ nd=0.00000E+000    	lnd=0.00000E+000    	wnd=0.00000E+000
+ rsh=2.1    cj=9.34e-04    cjsw=2.41e-10    js=1e-08    pb=0.90
+ pbsw=0.90    mj=0.491    mjsw=0.222    wdf=0    dell=0

.END
